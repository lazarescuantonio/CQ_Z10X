module char_rom(
   input  logic   [7:0] addr,
   output logic [127:0] data
   );

   always_comb
      case(addr)
         default: data = 128'b0;

 // code x41 (A)
         8'h41: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b00010000;   //   *
         data[ 31: 24] = 8'b00111000;   //  ***
         data[ 39: 32] = 8'b01101100;   // ** **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11111110;   //*******
         data[ 71: 64] = 8'b11111110;   //*******
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11000110;   //**   **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x42 (B)
         8'h42: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8]= 8'b00000000;   //
         data[ 23: 16]= 8'b11111100;   //******
         data[ 31: 24]= 8'b11111110;   //*******
         data[ 39: 32]= 8'b11000110;   //**   **
         data[ 47: 40]= 8'b11000110;   //**   **
         data[ 55: 48]= 8'b11111100;   //******
         data[ 63: 56]= 8'b11111100;   //******
         data[ 71: 64]= 8'b11000110;   //**   **
         data[ 79: 72]= 8'b11000110;   //**   **
         data[ 87: 80]= 8'b11111110;   //*******
         data[ 95: 88]= 8'b11111100;   //******
         data[103: 96]= 8'b00000000;   //
         data[111:104]= 8'b00000000;   //
         data[119:112]= 8'b00000000;   //
         data[127:120]= 8'b00000000;   //
         end
 // code x43 (C)
         8'h43: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b01111100;   // *****
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000000;   //**
         data[ 47: 40] = 8'b11000000;   //**
         data[ 55: 48] = 8'b11000000;   //**
         data[ 63: 56] = 8'b11000000;   //**
         data[ 71: 64] = 8'b11000000;   //**
         data[ 79: 72] = 8'b11000000;   //**
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b01111100;   // *****
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x44 (D)
         8'h44: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111100;   //******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b11111100;   //******
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x45 (E)
         8'h45: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000000;   //**
         data[ 47: 40] = 8'b11000000;   //**
         data[ 55: 48] = 8'b11111100;   //******
         data[ 63: 56] = 8'b11111100;   //******
         data[ 71: 64] = 8'b11000000;   //**
         data[ 79: 72] = 8'b11000000;   //**
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b11111110;   //*******
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x46 (F)
         8'h46: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000000;   //**
         data[ 47: 40] = 8'b11000000;   //**   
         data[ 55: 48] = 8'b11111100;   //******
         data[ 63: 56] = 8'b11111100;   //******
         data[ 71: 64] = 8'b11000000;   //** 
         data[ 79: 72] = 8'b11000000;   //** 
         data[ 87: 80] = 8'b11000000;   //**
         data[ 95: 88] = 8'b11000000;   //**
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x47 (G)
         8'h47: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b01111100;   // *****
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000000;   //**
         data[ 47: 40] = 8'b11000000;   //**   
         data[ 55: 48] = 8'b11111110;   //*******
         data[ 63: 56] = 8'b11111110;   //*******
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b01110110;   // *** **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x48 (H)
         8'h48: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11111110;   //*******
         data[ 63: 56] = 8'b11111110;   //*******
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11000110;   //**   **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x49 (I)
         8'h49: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b00110000;   //  **
         data[ 47: 40] = 8'b00110000;   //  **
         data[ 55: 48] = 8'b00110000;   //  **
         data[ 63: 56] = 8'b00110000;   //  **
         data[ 71: 64] = 8'b00110000;   //  **
         data[ 79: 72] = 8'b00110000;   //  **
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b11111110;   //*******
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4a (J)
         8'h4a: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b00011000;   //   **
         data[ 47: 40] = 8'b00011000;   //   **
         data[ 55: 48] = 8'b00011000;   //   **
         data[ 63: 56] = 8'b00011000;   //   **
         data[ 71: 64] = 8'b00011000;   //   **
         data[ 79: 72] = 8'b00011000;   //   **
         data[ 87: 80] = 8'b11111000;   //*****
         data[ 95: 88] = 8'b01111000;   // ****
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4b (K)
         8'h4b: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11001100;   //**  **
         data[ 39: 32] = 8'b11011000;   //** **
         data[ 47: 40] = 8'b11110000;   //****
         data[ 55: 48] = 8'b11100000;   //***
         data[ 63: 56] = 8'b11100000;   //***
         data[ 71: 64] = 8'b11110000;   //****
         data[ 79: 72] = 8'b11011000;   //** **
         data[ 87: 80] = 8'b11001100;   //**  **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4c (L)
         8'h4c: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000000;   //**
         data[ 31: 24] = 8'b11000000;   //**
         data[ 39: 32] = 8'b11000000;   //**
         data[ 47: 40] = 8'b11000000;   //**
         data[ 55: 48] = 8'b11000000;   //**
         data[ 63: 56] = 8'b11000000;   //**
         data[ 71: 64] = 8'b11000000;   //**
         data[ 79: 72] = 8'b11000000;   //**
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b11111110;   //*******
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4d (M)
         8'h4d: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11101110;   //*** ***
         data[ 47: 40] = 8'b11111110;   //*******
         data[ 55: 48] = 8'b11010110;   //** * **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11000110;   //**   **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4e (N)
         8'h4e: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11100110;   //***  **
         data[ 47: 40] = 8'b11110110;   //**** **
         data[ 55: 48] = 8'b11111110;   //*******
         data[ 63: 56] = 8'b11011110;   //** ****
         data[ 71: 64] = 8'b11001110;   //**  ***
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11000110;   //**   **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x4f (O)
         8'h4f: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b01111100;   // *****
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b01111100;   // *****
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x50 (P)
         8'h50: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111100;   //******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11111110;   //*******
         data[ 63: 56] = 8'b11111100;   //******   
         data[ 71: 64] = 8'b11000000;   //**   
         data[ 79: 72] = 8'b11000000;   //**   
         data[ 87: 80] = 8'b11000000;   //**
         data[ 95: 88] = 8'b11000000;   //**
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x51 (Q)
         8'h51: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111100;   // *****
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **  
         data[ 71: 64] = 8'b11010110;   //** * **
         data[ 79: 72] = 8'b11111110;   //*******
         data[ 87: 80] = 8'b01101100;   // ** ** 
         data[ 95: 88] = 8'b00000110;   //     **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x52 (R)
         8'h52: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111100;   //******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11111110;   //*******
         data[ 63: 56] = 8'b11111100;   //******   
         data[ 71: 64] = 8'b11011000;   //** **  
         data[ 79: 72] = 8'b11001100;   //**  ** 
         data[ 87: 80] = 8'b11000110;   //**   **
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x53 (S)
         8'h53: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b01111100;   // *****
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b11000000;   //**   
         data[ 47: 40] = 8'b11000000;   //**   
         data[ 55: 48] = 8'b11111100;   //******
         data[ 63: 56] = 8'b01111110;   // ******   
         data[ 71: 64] = 8'b00000110;   //     **  
         data[ 79: 72] = 8'b00000110;   //     **
         data[ 87: 80] = 8'b11111110;   //*******  
         data[ 95: 88] = 8'b01111100;   // ***** 
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x54 (T)
         8'h54: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b00110000;   //  **
         data[ 47: 40] = 8'b00110000;   //  **
         data[ 55: 48] = 8'b00110000;   //  **
         data[ 63: 56] = 8'b00110000;   //  **   
         data[ 71: 64] = 8'b00110000;   //  **  
         data[ 79: 72] = 8'b00110000;   //  **
         data[ 87: 80] = 8'b00110000;   //  **  
         data[ 95: 88] = 8'b00110000;   //  **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x55 (U)
         8'h55: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b11000110;   //**   **
         data[ 87: 80] = 8'b11111110;   //*******
         data[ 95: 88] = 8'b01111100;   // *****
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x56 (V)
         8'h56: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11000110;   //**   **
         data[ 79: 72] = 8'b01101100;   // ** **
         data[ 87: 80] = 8'b00111000;   //  ***  
         data[ 95: 88] = 8'b00010000;   //   * 
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x57 (W)
         8'h57: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b11000110;   //**   **
         data[ 47: 40] = 8'b11000110;   //**   **
         data[ 55: 48] = 8'b11000110;   //**   **
         data[ 63: 56] = 8'b11000110;   //**   **
         data[ 71: 64] = 8'b11010110;   //** * **
         data[ 79: 72] = 8'b11111110;   //*******
         data[ 87: 80] = 8'b11101110;   //*** ***  
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x58 (X)
         8'h58: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b01101100;   // ** ** 
         data[ 47: 40] = 8'b00111000;   //  ***
         data[ 55: 48] = 8'b00111000;   //  *** 
         data[ 63: 56] = 8'b00111000;   //  ***
         data[ 71: 64] = 8'b00111000;   //  ***
         data[ 79: 72] = 8'b01101100;   // ** **
         data[ 87: 80] = 8'b11000110;   //**   **  
         data[ 95: 88] = 8'b11000110;   //**   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x59 (Y)
         8'h59: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11000110;   //**   **
         data[ 31: 24] = 8'b11000110;   //**   **
         data[ 39: 32] = 8'b01101100;   // ** ** 
         data[ 47: 40] = 8'b00111000;   //  ***
         data[ 55: 48] = 8'b00011000;   //   ** 
         data[ 63: 56] = 8'b00011000;   //   **
         data[ 71: 64] = 8'b00011000;   //   **
         data[ 79: 72] = 8'b00011000;   //   **
         data[ 87: 80] = 8'b00011000;   //   **  
         data[ 95: 88] = 8'b00011000;   //   **
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
 // code x5a (Z)
         8'h5a: begin
         data[  7:  0] = 8'b00000000;   //
         data[ 15:  8] = 8'b00000000;   //
         data[ 23: 16] = 8'b11111110;   //*******
         data[ 31: 24] = 8'b11111110;   //*******
         data[ 39: 32] = 8'b00000110;   //     **  
         data[ 47: 40] = 8'b00001100;   //    **
         data[ 55: 48] = 8'b00011000;   //   ** 
         data[ 63: 56] = 8'b00110000;   //  **
         data[ 71: 64] = 8'b01100000;   // **
         data[ 79: 72] = 8'b11000000;   //**
         data[ 87: 80] = 8'b11111110;   //*******  
         data[ 95: 88] = 8'b11111110;   //*******
         data[103: 96] = 8'b00000000;   //
         data[111:104] = 8'b00000000;   //
         data[119:112] = 8'b00000000;   //
         data[127:120] = 8'b00000000;   //
         end
         
      endcase
endmodule